`define CLK_CYCLE      10000 
//`define CLK_CYCLE      0.9 
`define SETUP_CYCLE    0.1
`define RESET_CYCLE    18.3
